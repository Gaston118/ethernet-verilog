module shiftreg (
    output [3:0] o_led,
    input i_valid,
    input rst, 
    input clk
);

endmodule