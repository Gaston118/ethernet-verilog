module count (
    output o_valid,
    input [2:0] i_sw,
    input rst,
    input clk
);

endmodule